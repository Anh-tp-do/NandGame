module v_nand


endmdule

//

module v_invert 

endmodule

module v_and 

endmodule

module v_or 

endmodule

module v_xor 

endmodule
